module top_test_tb;

reg [3:0] a4bit,
reg  a16bit;
reg  clock, enable;
reg  q4bit;
reg q16bit;
    
endmodule