module c_addsub_0 (
  input [7:0] A,
  input [7:0] B,
  output wire [7:0] S
);
  
endmodule

module c_addsub_1 (
  input [7:0] A,
  input [7:0] B,
  output wire [7:0] S
);
  
endmodule

module c_addsub_2 (
  input [7:0] A,
  input [7:0] B,
  output wire [7:0] S
);
  
endmodule